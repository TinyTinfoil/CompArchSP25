`define CODE "code/blink.txt"
