`define CODE "code/code.txt"
